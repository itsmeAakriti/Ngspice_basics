* Netlist 

.include TSMC_180nm.txt
.param SUPPLY=1.8V
.param LAMBDA=0.09u
.param width_N=1.8u
.global gnd vdd

Vin a gnd pulse(0 1.8 0ns 100ps 100ps 9.9ns 20ns)
Vds vdd 0 'SUPPLY'
Cl c gnd 100fF

MP1 b a vdd gnd CMOSP W={2.5*width_N} L={4*LAMBDA} AS={5*width_N*LAMBDA} 
+ PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
MN1 b a gnd gnd CMOSN W={width_N} L={4*LAMBDA} AS={5*width_N*LAMBDA} 
+ PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

MP2 c b vdd gnd CMOSP W={2.5*width_N} L={4*LAMBDA} AS={5*width_N*LAMBDA} 
+ PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
MN2 c b gnd gnd CMOSN W={width_N} L={4*LAMBDA} AS={5*width_N*LAMBDA} 
+ PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

.tran 20n 40n 
.measure tran t_rise 
+TRIG AT=0.05n TARG v(C) VAL=0.7 RISE=1 CROSS=1
.measure tran t_fall 
+TRIG AT=10n TARG v(C) VAL=0.7 FALL=1 CROSS=2
.control  
run
set color0=white
set color1=black
plot v(c) v(a)

.endc
